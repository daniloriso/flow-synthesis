--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DYNAMIC_ADD_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT (
		CLOCK    :IN  STD_LOGIC;
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_ADD_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
  INPUT_2p  : STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		OUTPUT <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_1p),OUTPUT_1_WIDTH) - RESIZE(SIGNED(INPUT_2p),OUTPUT_1_WIDTH) );
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		OUTPUT <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_1p),OUTPUT_1_WIDTH) - RESIZE(SIGNED(INPUT_2p),OUTPUT_1_WIDTH) );
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  SUBSTRACTOR COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DYNAMIC_SUB_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		CLOCK    :IN  STD_LOGIC;
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_SUB_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
  INPUT_2p  : STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		OUTPUT <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1p),OUTPUT_1_WIDTH) - RESIZE(UNSIGNED(INPUT_2p),OUTPUT_1_WIDTH) );
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		OUTPUT <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_1p),OUTPUT_1_WIDTH) - RESIZE(SIGNED(INPUT_2p),OUTPUT_1_WIDTH) );
      END IF; -- IF(clock...)
      OUTPUT_1 <= OUTPUT_1p;
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DYNAMIC_MUL_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		CLOCK    :IN  STD_LOGIC;
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_MUL_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
  INPUT_2p  : STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
        OUTPUT <= STD_LOGIC_VECTOR(RESIZE(UNSIGNED(INPUT_1p) * UNSIGNED(INPUT_2p), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
        OUTPUT <= STD_LOGIC_VECTOR(RESIZE(SIGNED(INPUT_1p) * SIGNED(INPUT_2p), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#
--#
--#
--#
--####################################################################################################

--	MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DIVIDER_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DIVIDER_Dynamic IS
  -- MAXIMUM FUNCTION TO COMPUTE THE INTERNAL DATA SIZE
  FUNCTION maximum (left, right : NATURAL) return NATURAL IS
  BEGIN  -- function max
    IF LEFT > RIGHT THEN RETURN LEFT;
    ELSE RETURN RIGHT;
    END IF;
  END FUNCTION maximum;

BEGIN
	PROCESS (INPUT_1, INPUT_2)
		VARIABLE Stmp  : SIGNED  ((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
	begin
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED( INPUT_1 ) * UNSIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		ELSE
			Stmp     := RESIZE( SIGNED( INPUT_1 ) * SIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		END IF;
	END PROCESS;
END;


--####################################################################################################
--#
--#  MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;


ENTITY DYNAMIC_SQR_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		CLOCK    :IN  STD_LOGIC;
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_SQR_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        OUTPUT_1 <= STD_LOGIC_VECTOR(RESIZE(UNSIGNED(INPUT_1p) * UNSIGNED(INPUT_1p), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        OUTPUT_1 <= STD_LOGIC_VECTOR(RESIZE(SIGNED(INPUT_1p) * SIGNED(INPUT_1p), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#
--#
--#
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DYNAMIC_ABS_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_ABS_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        OUTPUT_1 <= STD_LOGIC_VECTOR(RESIZE( UNSIGNED(INPUT_1), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        OUTPUT_1 <= STD_LOGIC_VECTOR(RESIZE( abs(SIGNED( INPUT_1p)), OUTPUT_1_WIDTH));
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#
--#
--#
--#
--####################################################################################################

LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY RSHIFT_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF RSHIFT_Dynamic IS
BEGIN
	PROCESS (INPUT_1, INPUT_2)
		VARIABLE Stmp  : SIGNED  ((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
	begin
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED( INPUT_1 ) * UNSIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		ELSE
			Stmp     := RESIZE( SIGNED( INPUT_1 ) * SIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		END IF;
	END PROCESS;
END;


--####################################################################################################
--#
--#
--#
--#
--#
--####################################################################################################
--	MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY DYNAMIC_MAX_PIPELINE IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF DYNAMIC_MAX_PIPELINE IS
  INPUT_1p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
  INPUT_2p  : STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
BEGIN
	USIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		IF( UNSIGNED(INPUT_1p) > UNSIGNED(INPUT_2p) ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1p), OUTPUT_1_WIDTH) );
		ELSE
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_2p), OUTPUT_1_WIDTH) );
		END IF;
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (CLOCK)
	BEGIN
      IF ( clock'event AND clock = '1' ) THEN
        INPUT_1p  <= INPUT_1;
        INPUT_2p  <= INPUT_2;
		IF( SIGNED(INPUT_1p) > SIGNED(INPUT_2p) ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_1p), OUTPUT_1_WIDTH) );
		ELSE
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_2p), OUTPUT_1_WIDTH) );
		END IF;
      END IF; -- IF(clock...)
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#
--#
--#
--#
--####################################################################################################

--	MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY MIN_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF MIN_Dynamic IS
BEGIN
	USIG: IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		IF( UNSIGNED(INPUT_1) < UNSIGNED(INPUT_2) ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1), OUTPUT_1_WIDTH) );
		ELSE
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_2), OUTPUT_1_WIDTH) );
		END IF;
	END PROCESS;
	END GENERATE USIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		IF( SIGNED(INPUT_1) < SIGNED(INPUT_2) ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_1), OUTPUT_1_WIDTH) );
		ELSE
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(SIGNED(INPUT_2), OUTPUT_1_WIDTH) );
		END IF;
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY AND_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF AND_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) AND UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( SIGNED( INPUT_1 ) AND SIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY NAND_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF NAND_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) NAND UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( SIGNED( INPUT_1 ) NAND SIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY OR_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF OR_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) OR UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( SIGNED( INPUT_1 ) OR SIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY NOR_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF OR_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) NOR UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( SIGNED( INPUT_1 ) NOR SIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY XOR_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF XOR_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) XOR UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( SIGNED( INPUT_1 ) XOR SIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY NOT_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF XOR_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( NOT RESIZE( UNSIGNED( INPUT_1 ), OUTPUT_1_WIDTH ) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( NOT RESIZE( UNSIGNED( INPUT_1 ), OUTPUT_1_WIDTH ) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY absADD_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF absADD_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) + UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( ABS(SIGNED( INPUT_1 ) + SIGNED( INPUT_2 )), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;

--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY absSUB_Dynamic IS
  GENERIC(
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF absSUB_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) - UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( ABS(SIGNED( INPUT_1 ) - SIGNED( INPUT_2 )), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;


--####################################################################################################
--#
--#  ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--#  DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--#	 IMS LABORATORY -  UMR-CNRS 5218
--#
--####################################################################################################
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY rSHIFT_Dynamic IS
  GENERIC(
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF rSHIFT_Dynamic IS
BEGIN
	SIG:  IF C_SIGNED = 0 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		IF( UNSIGNED(INPUT_2) == 0 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 1 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 1)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 2 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 2)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 3 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 3)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 4 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 4)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 5 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 5)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 6 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 6)), OUTPUT_1_WIDTH) );
		ELSIF( UNSIGNED(INPUT_2) == 7 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 7)), OUTPUT_1_WIDTH) );
SIZE8:  IF INPUT_1'LENGTH > 8 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 8 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 8)), OUTPUT_1_WIDTH) );
END GENERATE SIZE8;
SIZE9:  IF INPUT_1'LENGTH > 9 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 9 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 9)), OUTPUT_1_WIDTH) );
END GENERATE SIZE9;
SIZE10: IF INPUT_1'LENGTH > 10 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 10 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 10)), OUTPUT_1_WIDTH) );
END GENERATE SIZE10;
SIZE11: IF INPUT_1'LENGTH > 11 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 11 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 11)), OUTPUT_1_WIDTH) );
END GENERATE SIZE11;
SIZE12: IF INPUT_1'LENGTH > 12 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 12 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 12)), OUTPUT_1_WIDTH) );
END GENERATE SIZE12;
SIZE13: IF INPUT_1'LENGTH > 13 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 13 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 13)), OUTPUT_1_WIDTH) );
END GENERATE SIZE13;
SIZE14: IF INPUT_1'LENGTH > 14 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 14 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 14)), OUTPUT_1_WIDTH) );
END GENERATE SIZE14;
SIZE15: IF INPUT_1'LENGTH > 15 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 15 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 15)), OUTPUT_1_WIDTH) );
END GENERATE SIZE15;
SIZE16: IF INPUT_1'LENGTH > 16 GENERATE
		ELSIF( UNSIGNED(INPUT_2) == 16 ) THEN
			OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE(UNSIGNED(INPUT_1(INPUT_1_WIDTH-1 DOWNTO 16)), OUTPUT_1_WIDTH) );
END GENERATE SIZE16;
		ELSE
			ASSERT (UNSIGNED(INPUT_2) == 16) FATAL "UN-MANAGED CASE IN THE RIGHT SHIFT OPERATOR";
		END IF;
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( UNSIGNED( INPUT_1 ) - UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;

	SIG:  IF C_SIGNED = 1 GENERATE
	PROCESS (INPUT_1, INPUT_2)
	BEGIN
		OUTPUT_1 <= STD_LOGIC_VECTOR( RESIZE( ABS(SIGNED( INPUT_1 ) - SIGNED( INPUT_2 )), OUTPUT_1_WIDTH) );
	END PROCESS;
	END GENERATE SIG;
END;
